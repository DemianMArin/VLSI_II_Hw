module mux32(
  input logic [31:0] a,
  input logic [31:0] b,
  input logic sel,
  output logic [31:0] y
);

endmodule
