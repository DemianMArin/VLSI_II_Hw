module Pri_En(
  input logic [7:0] D,
  output logic [2:0] Q
);

endmodule
